# ====================================================================
#
#      hal_arm_arm9_smdk2440.cdl
#
#      Samsung ARM9/smdk2440 evaluation board HAL package configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      michael anburaj <michaelanburaj@hotmail.com>
# Contributors:   michael anburaj <michaelanburaj@hotmail.com>
# Date:           2003-08-01
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_ARM_ARM9_SMDK2440 {
    display       "Samsung ARM9/smdk2440 development board"
    parent        CYGPKG_HAL_ARM_ARM9
    requires      CYGPKG_HAL_ARM_ARM9_ARM920T
    hardware
    include_dir   cyg/hal
    define_header hal_arm_arm9_smdk2440.h
    description   "
         The smdk2440 HAL package provides the support needed to run eCos on Samsung
         S3C2440X (ARM920T) based boards."

    compile       smdk2440_misc.c hal_diag.c

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    implements    CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_arm.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_VARIANT_H  <pkgconf/hal_arm_arm9.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_arm_arm9_smdk2440.h>"
        puts $::cdl_header "#define HAL_PLATFORM_CPU    \"ARM9\""
        puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"smdk2440 system\""
        puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"\""

        puts $::cdl_header "#define HAL_PLATFORM_MACHINE_TYPE  106"
    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        legal_values  { "RAM" "ROM" "ROMRAM" }
        default_value  { "ROM" }
        no_define
        define -file system.h CYG_HAL_STARTUP
        description   "
            When targetting the smdk2440 evaluation board it is possible to build
            the system for either RAM bootstrap or ROM bootstrap(s). Select
            'ram' when building programs to load into RAM using eCos GDB stubs.
            Select 'rom' when building a stand-alone application which will be
            put into ROM, or for the special case of building the eCos GDB stubs
            themselves."
    }

    # Both PLLs are in bypass mode on startup.
    # FIXME: Add proper configury
    cdl_option CYGNUM_HAL_ARM_SMDK2440_CPU_CLOCK {
        display       "CPU speed"
        flavor        data
        legal_values  176000000 180000000 184000000 192000000 200000000 405000000
        default_value { 405000000 }
        description   "
            This is the actual CPU operating frequency (FCLK)."
    }

    cdl_option CYGNUM_HAL_ARM_SMDK2440_BUS_CLOCK {
        display       "ARM920T bus speed"
        flavor        data
        calculated    { CYGNUM_HAL_ARM_SMDK2440_CPU_CLOCK / 3 }
        description   "
            This is the ARM920T AHB bus operating frequency (HCLK)."
    }

    cdl_option CYGNUM_HAL_ARM_SMDK2440_PERIPHERAL_CLOCK {
        display       "Peripheral bus speed"
        flavor        data
        calculated    { CYGNUM_HAL_ARM_SMDK2440_CPU_CLOCK / 6 }
        description   "
            This is the peripheral (APB) bus operating frequency (PCLK)."
    }

    cdl_option CYGNUM_HAL_ARM_SMDK2440_TIMER_PRESCALE {
        display       "Timer prescale"
        flavor        data
        legal_values  0 to 255
        default_value 16
        description   "
            This is the prescale value used on the clock used to drive
            the kernel counter. Note that some parts of the code may fail
            if this is changed due to over/underflows of expressions."
    }

    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants"
        flavor        none
        no_define
    
        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            calculated    1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            calculated    100
        }
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
            calculated    ((CYGNUM_HAL_ARM_SMDK2440_PERIPHERAL_CLOCK/CYGNUM_HAL_ARM_SMDK2440_TIMER_PRESCALE/2)/CYGNUM_HAL_RTC_DENOMINATOR)
            description   "
            Assuming 1/2 post prescale divider."
        }
    }

    cdl_component CYGSEM_SMDK2440_LCD_SUPPORT {
        display        "Support LCD"
        flavor         bool
        default_value  1
        compile        lcd_support.c
        description    "
          Enabling this option will enable the use the LCD as a 
          simple framebuffer, suitable for use with a windowing
          package."

    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD {
        display       "Diagnostic serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200
        default_value 115200
        description   "
            This option selects the baud rate used for the diagnostic port.
            Note: this should match the value chosen for the GDB port if the
            diagnostic and GDB port are the same."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_BAUD {
        display       "GDB serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200
        default_value 115200
        description   "
            This option selects the baud rate used for the diagnostic port.
            Note: this should match the value chosen for the GDB port if the
            diagnostic and GDB port are the same."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display      "Number of communication channels on the board"
        flavor       data
        calculated   2
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_DEFAULT {
        display      "Default console channel."
        flavor       data
        legal_values 0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        calculated   0
    }
 
    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_CONFIGURABLE
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
            The smdk2440 boards have two serial ports. This option
            chooses which port will be used to connect to a host
            running GDB."
     }
 
     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
         display         "Diagnostic serial port"
         active_if       CYGPRI_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_CONFIGURABLE
         flavor data
         legal_values    0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
         default_value   CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_DEFAULT
         description     "
             The smdk2440 boards have two serial ports.  This option
             chooses which port will be used for diagnostic output."
     }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        no_define
        description   "
            Global build options including control over
            compiler flags, linker flags and choice of toolchain."

        parent  CYGPKG_NONE

        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "arm-elf" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { "-mcpu=arm9 -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" }
            description   "
                This option controls the global compiler flags which are used to
                compile all packages by default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { "--no-target-default-spec -Wl,--gc-sections -Wl,-static -g -O2 -nostdlib" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }

        cdl_option CYGBLD_BUILD_GDB_STUBS {
            display "Build GDB stub ROM image"
            default_value 0
            requires { CYG_HAL_STARTUP == "ROM" }
            requires CYGSEM_HAL_ROM_MONITOR
            requires CYGBLD_BUILD_COMMON_GDB_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
            requires CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
            requires ! CYGDBG_HAL_COMMON_INTERRUPTS_SAVE_MINIMUM_CONTEXT
            requires ! CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM
            no_define
            description "
                This option enables the building of the GDB stubs for the
                board. The common HAL controls takes care of most of the
                build process, but the final conversion from ELF image to
                binary data is handled by the platform CDL, allowing
                relocation of the data if necessary."

            make -priority 320 {
                <PREFIX>/bin/gdb_module.bin : <PREFIX>/bin/gdb_module.img
                $(OBJCOPY) -O binary $< $@
            }
        }
   }


    cdl_component CYGPKG_HAL_ARM_ARM9_SMDK2440_OPTIONS {
        display "ARM9/smdk2440 build options"
        flavor  none
        no_define
        description   "
            Package specific build options including control over
            compiler flags used only in building this package,
            and details of which tests are built."

        cdl_option CYGPKG_HAL_ARM_ARM9_SMDK2440_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the ARM9 smdk2440 HAL. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_HAL_ARM_ARM9_SMDK2440_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the ARM9 smdk2440 HAL. These flags are removed from
                the set of global flags if present."
        }

        cdl_option CYGPKG_HAL_ARM_ARM9_SMDK2440_TESTS {
            display "ARM9/smdk2440 tests"
            flavor  data
            no_define
            calculated { "" }
            description   "
                This option specifies the set of tests for the ARM9/smdk2440 HAL."
        }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { CYG_HAL_STARTUP == "RAM" ? "arm_arm9_smdk2440_ram" : \
                     CYG_HAL_STARTUP == "ROM" ? "arm_arm9_smdk2440_rom" : \
                                                "arm_arm9_smdk2440_romram" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated {CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_arm9_smdk2440_ram.ldi>" :  \
                        CYG_HAL_STARTUP == "ROM" ? "<pkgconf/mlt_arm_arm9_smdk2440_rom.ldi>" : \
                                                   "<pkgconf/mlt_arm_arm9_smdk2440_romram.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_arm9_smdk2440_ram.h>" :  \
                         CYG_HAL_STARTUP == "ROM" ? "<pkgconf/mlt_arm_arm9_smdk2440_rom.h>" : \
                                                    "<pkgconf/mlt_arm_arm9_smdk2440_romram.h>" }
        }
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { (CYG_HAL_STARTUP == "ROM") || (CYG_HAL_STARTUP == "ROMRAM") }
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }

    cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
         display       "Work with a ROM monitor"
         flavor        booldata
         legal_values  { "GDB_stubs" }
         default_value { CYG_HAL_STARTUP == "RAM" ? "GDB_stubs" : 0 }
         parent        CYGPKG_HAL_ROM_MONITOR
         requires      { CYG_HAL_STARTUP == "RAM" }
         description   "
             Support can be enabled for different varieties of ROM monitor.
             This support changes various eCos semantics such as the encoding
             of diagnostic output, or the overriding of hardware interrupt
             vectors.
             \"GDB_stubs\" provides support when GDB stubs are included in
             the ROM monitor or boot ROM."
     }

    cdl_component CYGPKG_REDBOOT_HAL_OPTIONS {
        display       "Redboot HAL options"
        flavor        none
        no_define
        parent        CYGPKG_REDBOOT
        active_if     CYGPKG_REDBOOT
        description   "
            This option lists the target's requirements for a valid Redboot
            configuration."

        # The backup image is not needed, since ROMRAM is the normal
        # RedBoot startup type.
        requires {!CYGPKG_REDBOOT_FLASH || CYGOPT_REDBOOT_FIS_REDBOOT_BACKUP == 0}

        # RedBoot details
        requires { CYGPKG_REDBOOT_ARM_LINUX_EXEC }
        requires { CYGHWR_REDBOOT_ARM_LINUX_EXEC_ADDRESS_DEFAULT == 0x00008000 }
        define_proc {
            puts $::cdl_header "#define CYGHWR_REDBOOT_ARM_TRAMPOLINE_ADDRESS 0x00001f00"
        }
    
        cdl_option CYGBLD_BUILD_REDBOOT_BIN {
            display       "Build Redboot ROM binary image"
            active_if     CYGBLD_BUILD_REDBOOT
            default_value 1
            no_define
            description "This option enables the conversion of the Redboot ELF
                         image to a binary image suitable for ROM programming."
    
            make -priority 325 {
                <PREFIX>/bin/redboot.bin : <PREFIX>/bin/redboot.elf
                $(OBJCOPY) --strip-debug $< $(@:.bin=.img) 
                $(OBJCOPY) -O srec $< $(@:.bin=.srec)
                $(OBJCOPY) -O binary $< $@
            }
        }
    }

}
 